module REG_FILE_tb;

endmodule
