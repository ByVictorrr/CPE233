`include "./RAT_MCU.sv"
/*
 * RAT_MCU_tb
 * Copyright (C) 2019 victor <victor@TheShell>
 *
 * Distributed under terms of the MIT license.
 */

//////////////////////////////////////////////////////////////////////////////////
// Engineer: Victor Delaplaine
// 
// Create Date: 02/07/2019 20:38
// Design Name: 
// Module Name: RAT_MCU_tb
// Project Name: 
// Target Devices: Basy3 
// Tool Versions: 
// Description: 
// 		
// Dependencies: 
// 
// Revision:
// Revision 1.00 - File Created (02-07-2019) 
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RAT_MCU_tb();

	
	logic [7:0] IN_PORT;
	logic RESET;
	logic INT;
	logic CLK(CLK);
	logic [7:0] OUT_PORT;
	logic [7:0] PORT_ID;
	logic IO_STRB;



	RAT_MCU MCU( 
endmodule

