module SCTRACH_RAM_tb;

endmodule
